module pad_core_gnd();
// this is a wrapper
 VSS VSS_pad_local(GND,VDDIO,VDD,GNDIO);
  
endmodule // pad_core_gnd

module pad_core_vdd();
// this is a wrapper
VDD VDD_pad_local(GND,VDDIO,VDD,GNDIO);
   
endmodule // pad_vdd
